`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module transparent_d_latch (output logic q, input logic d, input logic c);

	// add code here
	lvl_sen_sr_latch u_lvl(.c,.r(~d),.s(d),.q);
endmodule
